CIRCUIT C:\users\huthayfa\Desktop\and.MSK
*
* IC Technology: CMOS 65nm general purpose - 8 Metal copper - strain - SiON oxide
*
VDD 1 0 DC 1.00
VB 7 0 DC 0 PULSE(0.00 1.00 0.04N 0.00N 0.00N 0.04N 0.08N)
VA 8 0 DC 0 PULSE(0.00 1.00 0.02N 0.00N 0.00N 0.02N 0.04N)
*
* List of nodes
* "A and B" corresponds to n�3
* "N4" corresponds to n�4
* "N6" corresponds to n�6
* "B" corresponds to n�7
* "A" corresponds to n�8
*
* MOS devices
MN1 0 4 3 0 N1  W= 0.35U L= 0.07U
MN2 6 8 0 0 N1  W= 0.38U L= 0.14U
MN3 4 7 6 0 N1  W= 0.35U L= 0.07U
MP1 1 4 3 1 P1  W= 0.49U L= 0.07U
MP2 4 8 1 1 P1  W= 0.49U L= 0.07U
MP3 1 7 4 1 P1  W= 0.52U L= 0.14U
*
C2 1 0  0.704fF
C3 3 0  0.294fF
C4 4 0  0.388fF
C6 6 0  0.105fF
C7 7 0  0.073fF
C8 8 0  0.122fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.35 U0=0.055 TOXE= 1.1E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.000
+DVT1=0.750 LPE0=0.200e-9 ETA0=0.080
+NFACTOR=  1.0 U0=0.055 UA=7.000e-15
+WINT=0.005U LPE0=0.200e-9 
+KT1=-0.050 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.32 U0=0.027 TOXE= 1.1E-9 LINT=0.010U 
+K1 =0.500 K2=0.100 DVT0=2.000
+DVT1=0.650 LPE0=0.200e-9 ETA0=0.080
+NFACTOR=  1.1 U0=0.027 UA=4.800e-15
+WINT=0.005U LPE0=0.200e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.010
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 1.00N
print  V(7) V(8) V(3) > out.txt
plot  V(7) V(8) V(3)
.endc
.END
